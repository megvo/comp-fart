//////////////////////////////////////////////////////////////////////////////////
// The Cooper Union
// ECE 251 Spring 2024
// Engineer: Megan Vo and Lamiah Khan
// 
//     Create Date: 2024-04-27
//     Module Name: datapath
//     Description: 32-bit RISC-based CPU datapath (MIPS)
//
// Revision: 1.0
//
//////////////////////////////////////////////////////////////////////////////////

`ifndef DATAPATH
`define DATAPATH

`timescale 1ns/100ps

`include "regfile.sv"
`include "alu.sv"
`include "dff.sv"
`include "adder.sv"
`include "sl2.sv"
`include "mux2.sv"
`include "signext.sv"

module datapath
    #(parameter n = 32)(
    //
    // ---------------- PORT DEFINITIONS ----------------
    //
    input  logic        clk, reset,
    input  logic [1:0]  memtoreg, 
    input  logic        pcsrc,
    input  logic        alusrc, 
    input  logic [1:0]  regdst, 
    input  logic        regwrite,
    input  logic [1:0]  jump,
    input  logic [2:0]  alucontrol,
    output logic        zero,
    output logic [(n-1):0] pc,
    input  logic [(n-1):0] instr,
    output logic [(n-1):0] aluout, writedata,
    input  logic [(n-1):0] readdata
);
    //
    // ---------------- MODULE DESIGN IMPLEMENTATION ----------------
    //
    logic [4:0]  writereg;
    logic [(n-1):0] pcnext, pcnextbr, pcplus4, pcbranch;
    logic [(n-1):0] signimm, signimmsh;
    logic [(n-1):0] srca, srcb;
    logic [(n-1):0] result;

    // "next PC" logic
    dff #(n)  pcreg(clk, reset, pcnext, pc);
  adder       pcadd1(.A(pc), .B(4), .Cin(1'b0), .Cout(Cout1), .Sum(pcplus4));
    sl2         immsh(signimm, signimmsh);
  adder       pcadd2(.A(pcplus4), .B(signimmsh), .Cin(1'b0), .Cout(Cout2), .Sum(pcbranch));
    mux2 #(n)   pcbrmux(pcplus4, pcbranch, pcsrc, pcnextbr);
    mux4 #(n)   pcmux(pcnextbr, {pcplus4[31:28], instr[25:0], 2'b00}, readdata, 32'hxxxxxxxx, jump, pcnext);

    // register file logic
    regfile     rf(clk, regwrite, instr[25:21], instr[20:16], writereg, result, srca, writedata);
    mux4 #(5)   wrmux(instr[20:16], instr[15:11], 5'b01111, 5'bxxxxx, regdst, writereg);
    mux4 #(n)   resmux(aluout, readdata, pcplus4, 32'hxxxxxxxx, memtoreg, result);
    signext     se(instr[15:0], signimm);

    // ALU logic
    mux2 #(n)   srcbmux(writedata, signimm, alusrc, srcb);
    alu         alu(clk, srca, srcb, alucontrol, aluout, zero);

endmodule

`endif // DATAPATH
